library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity I_CACHE is
    port(
        pc    : in  std_logic_vector(31 downto 0);
        instr : out std_logic_vector(31 downto 0)
    );
end I_CACHE;

architecture behavior of I_CACHE is
    signal address : std_logic_vector(4 downto 0);
begin

    address <= pc(4 downto 0);

    process(address)
    begin
        case address is

            ------------------------------------------------------------------
            -- 0: addi $1, $0, 5
            ------------------------------------------------------------------
            when "00000" =>  -- PC = 0
                instr <= "00100000000000010000000000000101";
                -- addi r1, r0, 5

            ------------------------------------------------------------------
            -- 1: addi $2, $0, 10
            ------------------------------------------------------------------
            when "00001" =>  -- PC = 1
                instr <= "00100000000000100000000000001010";
                -- addi r2, r0, 10

            ------------------------------------------------------------------
            -- 2: add $3, $1, $2   (r3 = 15)
            ------------------------------------------------------------------
            when "00010" =>  -- PC = 2
                instr <= "00000000001000100001100000100000";
                -- add r3, r1, r2

            ------------------------------------------------------------------
            -- 3: sub $4, $2, $1   (r4 = 5)
            ------------------------------------------------------------------
            when "00011" =>  -- PC = 3
                instr <= "00000000010000010010000000100010";
                -- sub r4, r2, r1

            ------------------------------------------------------------------
            -- 4: sw $3, 0($0)  (mem[0] = 15)
            ------------------------------------------------------------------
            when "00100" =>  -- PC = 4
                instr <= "10101100000000110000000000000000";
                -- sw r3, 0(r0)

            ------------------------------------------------------------------
            -- 5: lw $5, 0($0)  (r5 = 15, matches r3)
            ------------------------------------------------------------------
            when "00101" =>  -- PC = 5
                instr <= "10001100000001010000000000000000";
                -- lw r5, 0(r0)

            ------------------------------------------------------------------
            -- 6: init r6 = 0x2000_0000 (for overflow)
            ------------------------------------------------------------------
            when "00110" =>  -- PC = 6
                instr <= "00111100000001100010000000000000";
                -- lui r6, 0x2000   ; r6 = 0x20000000

            ------------------------------------------------------------------
            -- 7: r6 = r6 + r6  (Loop for overflow)
            ------------------------------------------------------------------
            when "00111" =>  -- PC = 7
                instr <= "00000000110001100011000000100000";
                -- add r6, r6, r6

            ------------------------------------------------------------------
            -- 8: beq r3, r5, +1  (15 == 15 → taken, skip PC9)
            ------------------------------------------------------------------
            when "01000" =>  -- PC = 8
                instr <= "00010000011001010000000000000001";
                -- beq r3, r5, +1

            ------------------------------------------------------------------
            -- 9: will be skipped if beq works
            ------------------------------------------------------------------
            when "01001" =>  -- PC = 9
                instr <= "00100000000001110000000000000001";
                -- addi r7, r0, 1   ; should be skipped

            ------------------------------------------------------------------
            -- 10: r7 = -1
            ------------------------------------------------------------------
            when "01010" =>  -- PC = 10
                instr <= "00100000000001111111111111111111";
                -- addi r7, r0, -1

            ------------------------------------------------------------------
            -- 11: bltz r7, +1 (taken, skip PC12)
            ------------------------------------------------------------------
            when "01011" =>  -- PC = 11
                instr <= "00000100111000000000000000000001";
                -- bltz r7, +1

            ------------------------------------------------------------------
            -- 12: skipped by bltz
            ------------------------------------------------------------------
            when "01100" =>  -- PC = 12
                instr <= "00100000000001100000000000101010";
                -- addi r6, r0, 42  ; should NOT execute

            ------------------------------------------------------------------
            -- 13: j 7 (loop back to overflow instruction)
            ------------------------------------------------------------------
            when "01101" =>  -- PC = 13
                instr <= "00001000000000000000000000000111";
                -- j 7

            ------------------------------------------------------------------
            -- Default: NOP
            ------------------------------------------------------------------
            when others =>
                instr <= (others => '0');  -- nop

        end case;
    end process;
end behavior;
